library ieee;
use ieee.std_logic_1164.all;

entity Exercise2 is
	port (a: in std_logic;
		b: in std_logic;
		o: out std_logic);
end entity;

architecture Behavioral of Exercise2 is
begin
	o <= ...;
end architecture;
